// Parameters for the Funct7 

`ifndef FUNCT7_PARAMETERS_VH
`define FUNCT7_PARAMETERS_VH

// Funct7 parameters
`define ADDFunct7 7'b0000000
`define SUBFunct7 7'b0100000
`define RS32MFunct7 7'b0000001
`define SetFunct7 7'b0000000
`define BitFunct7 7'b0000000
`define LogicalFunct7 7'b0000000
`define ArthematicFunct7 7'b0100000

`endif